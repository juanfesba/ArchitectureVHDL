LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity BCD is
port
(
	DataDer: in std_logic_vector(6 downto 0);
	DataIzq: in std_logic_vector(6 downto 0);
	SalidaData1: out std_logic_vector(6 downto 0);
	SalidaData2: out std_logic_vector(6 downto 0);
	SalidaData3: out std_logic_vector(6 downto 0);
	SalidaData4: out std_logic_vector(6 downto 0)
);
end entity;

architecture BCD of BCD is
begin
	process(DataDer, DataIzq)
		begin
			case DataDer is
			------- 0 al 9 -------------------
				when "0000000" => --0
					SalidaData1 <= "1000000"; --0
					SalidaData2 <= "1000000";
				when "0000001" => --1
					SalidaData1 <= "1111001"; --1
					SalidaData2 <= "1000000";
				when "0000010" => --2
					SalidaData1 <= "0100100"; --2
					SalidaData2 <= "1000000";
				when "0000011" => --3
					SalidaData1 <= "0110000"; --3
					SalidaData2 <= "1000000";
				when "0000100" => --4
					SalidaData1 <= "0011001"; --4
					SalidaData2 <= "1000000";
				when "0000101" => --5
					SalidaData1 <= "0010010"; --5
					SalidaData2 <= "1000000";
				when "0000110" => --6
					SalidaData1 <= "0000010"; --6
					SalidaData2 <= "1000000";
				when "0000111" => --7
					SalidaData1 <= "1111000"; --7
					SalidaData2 <= "1000000";
				when "0001000" => --8
					SalidaData1 <= "0000000"; --8
					SalidaData2 <= "1000000";
				when "0001001" => --9
					SalidaData1 <= "0010000"; --9
					SalidaData2 <= "1000000";
				------ 10 al 19 ----------------
				when "0001010" => --10
					SalidaData1 <= "1000000"; 
					SalidaData2 <= "1111001";
				when "0001011" => --11
					SalidaData1 <= "1111001";
					SalidaData2 <= "1111001";
				when "0001100" => --12
					SalidaData1 <= "0100100";
					SalidaData2 <= "1111001";
				when "0001101" => --13
					SalidaData1 <= "0110000";
					SalidaData2 <= "1111001";
				when "0001110" => --14
					SalidaData1 <= "0011001";
					SalidaData2 <= "1111001";
				when "0001111" => --15
					SalidaData1 <= "0010010";
					SalidaData2 <= "1111001";
				when "0010000" => --16
					SalidaData1 <= "0000010";
					SalidaData2 <= "1111001";
				when "0010001" => --17
					SalidaData1 <= "1111000";
					SalidaData2 <= "1111001";
				when "0010010" => --18
					SalidaData1 <= "0000000";
					SalidaData2 <= "1111001";
				when "0010011" => --19
					SalidaData1 <= "0010000";
					SalidaData2 <= "1111001";
				---- 20 al 29 -----------------
				when "0010100" => --20
					SalidaData1 <= "1000000";
					SalidaData2 <= "0100100";
				when "0010101" => --21
					SalidaData1 <= "1111001";
					SalidaData2 <= "0100100";
				when "0010110" => --22
					SalidaData1 <= "0100100";
					SalidaData2 <= "0100100";
				when "0010111" => --23
					SalidaData1 <= "0110000";
					SalidaData2 <= "0100100";
				when "0011000" => --24
					SalidaData1 <= "0011001";
					SalidaData2 <= "0100100";
				when "0011001" => --25
					SalidaData1 <= "0010010";
					SalidaData2 <= "0100100";
				when "0011010" => --26
					SalidaData1 <= "0000010";
					SalidaData2 <= "0100100";
				when "0011011" => --27
					SalidaData1 <= "1111000";
					SalidaData2 <= "0100100";
				when "0011100" => --28
					SalidaData1 <= "0000000";
					SalidaData2 <= "0100100";
				when "0011101" => --29
					SalidaData1 <= "0010000";
					SalidaData2 <= "0100100";
				---- 30 al 39 ----------------
				when "0011110" => --30
					SalidaData1 <= "1000000";
					SalidaData2 <= "0110000";
				when "0011111" => --31
					SalidaData1 <= "1111001";
					SalidaData2 <= "0110000";
				when "0100000" => --32
					SalidaData1 <= "0100100";
					SalidaData2 <= "0110000";
				when "0100001" => --33
					SalidaData1 <= "0110000";
					SalidaData2 <= "0110000";
				when "0100010" => --34
					SalidaData1 <= "0011001";
					SalidaData2 <= "0110000";
				when "0100011" => --35
					SalidaData1 <= "0010010";
					SalidaData2 <= "0110000";
				when "0100100" => --36
					SalidaData1 <= "0000010";
					SalidaData2 <= "0110000";
				when "0100101" => --37
					SalidaData1 <= "1111000";
					SalidaData2 <= "0110000";
				when "0100110" => --38
					SalidaData1 <= "0000000";
					SalidaData2 <= "0110000";
				when "0100111" => --39
					SalidaData1 <= "0010000";
					SalidaData2 <= "0110000";
				---- 40 al 49 --------------
				when "0101000" => --40
					SalidaData1 <= "1000000";
					SalidaData2 <= "0011001";
				when "0101001" => --41
					SalidaData1 <= "1111001";
					SalidaData2 <= "0011001";
				when "0101010" => --42
					SalidaData1 <= "0100100";
					SalidaData2 <= "0011001";
				when "0101011" => --43
					SalidaData1 <= "0110000";
					SalidaData2 <= "0011001";
				when "0101100" => --44
					SalidaData1 <= "0011001";
					SalidaData2 <= "0011001";
				when "0101101" => --45
					SalidaData1 <= "0010010";
					SalidaData2 <= "0011001";
				when "0101110" => --46
					SalidaData1 <= "0000010";
					SalidaData2 <= "0011001";
				when "0101111" => --47
					SalidaData1 <= "1111000";
					SalidaData2 <= "0011001";
				when "0110000" => --48
					SalidaData1 <= "0000000";
					SalidaData2 <= "0011001";
				when "0110001" => --49
					SalidaData1 <= "0010000";
					SalidaData2 <= "0011001";
				---- 50 al 59 ---------------
				when "0110010" => --50
					SalidaData1 <= "1000000";
					SalidaData2 <= "0010010";
				when "0110011" => --51
					SalidaData1 <= "1111001";
					SalidaData2 <= "0010010";
				when "0110100" => --52
					SalidaData1 <= "0100100";
					SalidaData2 <= "0010010";
				when "0110101" => --53
					SalidaData1 <= "0110000";
					SalidaData2 <= "0010010";
				when "0110110" => --54
					SalidaData1 <= "0011001";
					SalidaData2 <= "0010010";
				when "0110111" => --55
					SalidaData1 <= "0010010";
					SalidaData2 <= "0010010";
				when "0111000" => --56
					SalidaData1 <= "0000010";
					SalidaData2 <= "0010010";
				when "0111001" => --57
					SalidaData1 <= "1111000";
					SalidaData2 <= "0010010";
				when "0111010" => --58
					SalidaData1 <= "0000000";
					SalidaData2 <= "0010010";
				when "0111011" => --59
					SalidaData1 <= "0010000";
					SalidaData2 <= "0010010";
				---- 60 al 69 ---------------
				when "0111100" => --60
					SalidaData1 <= "1000000";
					SalidaData2 <= "0000010";
				when "0111101" => --61
					SalidaData1 <= "1111001";
					SalidaData2 <= "0000010";
				when "0111110" => --62
					SalidaData1 <= "0100100";
					SalidaData2 <= "0000010";
				when "0111111" => --63
					SalidaData1 <= "0110000";
					SalidaData2 <= "0000010";
				when "1000000" => --64
					SalidaData1 <= "0011001";
					SalidaData2 <= "0000010";
				when "1000001" => --65
					SalidaData1 <= "0010010";
					SalidaData2 <= "0000010";
				when "1000010" => --66
					SalidaData1 <= "0000010";
					SalidaData2 <= "0000010";
				when "1000011" => --67
					SalidaData1 <= "1111000";
					SalidaData2 <= "0000010";
				when "1000100" => --68
					SalidaData1 <= "0000000";
					SalidaData2 <= "0000010";
				when "1000101" => --69
					SalidaData1 <= "0010000";
					SalidaData2 <= "0000010";
				---- 70 al 79 ---------------
				when "1000110" => --70
					SalidaData1 <= "1000000";
					SalidaData2 <= "1111000";
				when "1000111" => --71
					SalidaData1 <= "1111001";
					SalidaData2 <= "1111000";
				when "1001000" => --72
					SalidaData1 <= "0100100";
					SalidaData2 <= "1111000";
				when "1001001" => --73
					SalidaData1 <= "0110000";
					SalidaData2 <= "1111000";
				when "1001010" => --74
					SalidaData1 <= "0011001";
					SalidaData2 <= "1111000";
				when "1001011" => --75
					SalidaData1 <= "0010010";
					SalidaData2 <= "1111000";
				when "1001100" => --76
					SalidaData1 <= "0000010";
					SalidaData2 <= "1111000";
				when "1001101" => --77
					SalidaData1 <= "1111000";
					SalidaData2 <= "1111000";
				when "1001110" => --78
					SalidaData1 <= "0000000";
					SalidaData2 <= "1111000";
				when "1001111" => --79
					SalidaData1 <= "0010000";
					SalidaData2 <= "1111000";
				---- 80 al 89 ---------------
				when "1010000" => --80
					SalidaData1 <= "1000000";
					SalidaData2 <= "0000000";
				when "1010001" => --81
					SalidaData1 <= "1111001";
					SalidaData2 <= "0000000";
				when "1010010" => --82
					SalidaData1 <= "0100100";
					SalidaData2 <= "0000000";
				when "1010011" => --83
					SalidaData1 <= "0110000";
					SalidaData2 <= "0000000";
				when "1010100" => --84
					SalidaData1 <= "0011001";
					SalidaData2 <= "0000000";
				when "1010101" => --85
					SalidaData1 <= "0010010";
					SalidaData2 <= "0000000";
				when "1010110" => --86
					SalidaData1 <= "0000010";
					SalidaData2 <= "0000000";
				when "1010111" => --87
					SalidaData1 <= "1111000";
					SalidaData2 <= "0000000";
				when "1011000" => --88
					SalidaData1 <= "0000000";
					SalidaData2 <= "0000000";
				when "1011001" => --89
					SalidaData1 <= "0010000";
					SalidaData2 <= "0000000";
				---- 80 al 89 ---------------
				when "1011010" => --90
					SalidaData1 <= "1000000";
					SalidaData2 <= "0010000";
				when "1011011" => --91
					SalidaData1 <= "1111001";
					SalidaData2 <= "0010000";
				when "1011100" => --92
					SalidaData1 <= "0100100";
					SalidaData2 <= "0010000";
				when "1011101" => --93
					SalidaData1 <= "0110000";
					SalidaData2 <= "0010000";
				when "1011110" => --94
					SalidaData1 <= "0011001";
					SalidaData2 <= "0010000";
				when "1011111" => --95
					SalidaData1 <= "0010010";
					SalidaData2 <= "0010000";
				when "1100000" => --96
					SalidaData1 <= "0000010";
					SalidaData2 <= "0010000";
				when "1100001" => --97
					SalidaData1 <= "1111000";
					SalidaData2 <= "0010000";
				when "1100010" => --98
					SalidaData1 <= "0000000";
					SalidaData2 <= "0010000";
				when "1100011" => --99
					SalidaData1 <= "0010000";
					SalidaData2 <= "0010000";
				when others =>
					SalidaData1 <= "1111111";
					SalidaData2 <= "1111111";
			end case;
			
			case DataIzq is
				when "0000000" => --0
					SalidaData3 <= "1000000"; --0
					SalidaData4 <= "1000000";
				when "0000001" => --1
					SalidaData3 <= "1111001"; --1
					SalidaData4 <= "1000000";
				when "0000010" => --2
					SalidaData3 <= "0100100"; --2
					SalidaData4 <= "1000000";
				when "0000011" => --3
					SalidaData3 <= "0110000"; --3
					SalidaData4 <= "1000000";
				when "0000100" => --4
					SalidaData3 <= "0011001"; --4
					SalidaData4 <= "1000000";
				when "0000101" => --5
					SalidaData3 <= "0010010"; --5
					SalidaData4 <= "1000000";
				when "0000110" => --6
					SalidaData3 <= "0000010"; --6
					SalidaData4 <= "1000000";
				when "0000111" => --7
					SalidaData3 <= "1111000"; --7
					SalidaData4 <= "1000000";
				when "0001000" => --8
					SalidaData3 <= "0000000"; --8
					SalidaData4 <= "1000000";
				when "0001001" => --9
					SalidaData3 <= "0010000"; --9
					SalidaData4 <= "1000000";
				------ 10 al 19 ----------------
				when "0001010" => --10
					SalidaData3 <= "1000000"; 
					SalidaData4 <= "1111001";
				when "0001011" => --11
					SalidaData3 <= "1111001";
					SalidaData4 <= "1111001";
				when "0001100" => --12
					SalidaData3 <= "0100100";
					SalidaData4 <= "1111001";
				when "0001101" => --13
					SalidaData3 <= "0110000";
					SalidaData4 <= "1111001";
				when "0001110" => --14
					SalidaData3 <= "0011001";
					SalidaData4 <= "1111001";
				when "0001111" => --15
					SalidaData3 <= "0010010";
					SalidaData4 <= "1111001";
				when "0010000" => --16
					SalidaData3 <= "0000010";
					SalidaData4 <= "1111001";
				when "0010001" => --17
					SalidaData3 <= "1111000";
					SalidaData4 <= "1111001";
				when "0010010" => --18
					SalidaData3 <= "0000000";
					SalidaData4 <= "1111001";
				when "0010011" => --19
					SalidaData3 <= "0010000";
					SalidaData4 <= "1111001";
				---- 20 al 29 -----------------
				when "0010100" => --20
					SalidaData3 <= "1000000";
					SalidaData4 <= "0100100";
				when "0010101" => --21
					SalidaData3 <= "1111001";
					SalidaData4 <= "0100100";
				when "0010110" => --22
					SalidaData3 <= "0100100";
					SalidaData4 <= "0100100";
				when "0010111" => --23
					SalidaData3 <= "0110000";
					SalidaData4 <= "0100100";
				when "0011000" => --24
					SalidaData3 <= "0011001";
					SalidaData4 <= "0100100";
				when "0011001" => --25
					SalidaData3 <= "0010010";
					SalidaData4 <= "0100100";
				when "0011010" => --26
					SalidaData3 <= "0000010";
					SalidaData4 <= "0100100";
				when "0011011" => --27
					SalidaData3 <= "1111000";
					SalidaData4 <= "0100100";
				when "0011100" => --28
					SalidaData3 <= "0000000";
					SalidaData4 <= "0100100";
				when "0011101" => --29
					SalidaData3 <= "0010000";
					SalidaData4 <= "0100100";
				---- 30 al 39 ----------------
				when "0011110" => --30
					SalidaData3 <= "1000000";
					SalidaData4 <= "0110000";
				when "0011111" => --31
					SalidaData3 <= "1111001";
					SalidaData4 <= "0110000";
				when "0100000" => --32
					SalidaData3 <= "0100100";
					SalidaData4 <= "0110000";
				when "0100001" => --33
					SalidaData3 <= "0110000";
					SalidaData4 <= "0110000";
				when "0100010" => --34
					SalidaData3 <= "0011001";
					SalidaData4 <= "0110000";
				when "0100011" => --35
					SalidaData3 <= "0010010";
					SalidaData4 <= "0110000";
				when "0100100" => --36
					SalidaData3 <= "0000010";
					SalidaData4 <= "0110000";
				when "0100101" => --37
					SalidaData3 <= "1111000";
					SalidaData4 <= "0110000";
				when "0100110" => --38
					SalidaData3 <= "0000000";
					SalidaData4 <= "0110000";
				when "0100111" => --39
					SalidaData3 <= "0010000";
					SalidaData4 <= "0110000";
				---- 40 al 49 --------------
				when "0101000" => --40
					SalidaData3 <= "1000000";
					SalidaData4 <= "0011001";
				when "0101001" => --41
					SalidaData3 <= "1111001";
					SalidaData4 <= "0011001";
				when "0101010" => --42
					SalidaData3 <= "0100100";
					SalidaData4 <= "0011001";
				when "0101011" => --43
					SalidaData3 <= "0110000";
					SalidaData4 <= "0011001";
				when "0101100" => --44
					SalidaData3 <= "0011001";
					SalidaData4 <= "0011001";
				when "0101101" => --45
					SalidaData3 <= "0010010";
					SalidaData4 <= "0011001";
				when "0101110" => --46
					SalidaData3 <= "0000010";
					SalidaData4 <= "0011001";
				when "0101111" => --47
					SalidaData3 <= "1111000";
					SalidaData4 <= "0011001";
				when "0110000" => --48
					SalidaData3 <= "0000000";
					SalidaData4 <= "0011001";
				when "0110001" => --49
					SalidaData3 <= "0010000";
					SalidaData4 <= "0011001";
				---- 50 al 59 ---------------
				when "0110010" => --50
					SalidaData3 <= "1000000";
					SalidaData4 <= "0010010";
				when "0110011" => --51
					SalidaData3 <= "1111001";
					SalidaData4 <= "0010010";
				when "0110100" => --52
					SalidaData3 <= "0100100";
					SalidaData4 <= "0010010";
				when "0110101" => --53
					SalidaData3 <= "0110000";
					SalidaData4 <= "0010010";
				when "0110110" => --54
					SalidaData3 <= "0011001";
					SalidaData4 <= "0010010";
				when "0110111" => --55
					SalidaData3 <= "0010010";
					SalidaData4 <= "0010010";
				when "0111000" => --56
					SalidaData3 <= "0000010";
					SalidaData4 <= "0010010";
				when "0111001" => --57
					SalidaData3 <= "1111000";
					SalidaData4 <= "0010010";
				when "0111010" => --58
					SalidaData3 <= "0000000";
					SalidaData4 <= "0010010";
				when "0111011" => --59
					SalidaData3 <= "0010000";
					SalidaData4 <= "0010010";
				---- 60 al 69 ---------------
				when "0111100" => --60
					SalidaData3 <= "1000000";
					SalidaData4 <= "0000010";
				when "0111101" => --61
					SalidaData3 <= "1111001";
					SalidaData4 <= "0000010";
				when "0111110" => --62
					SalidaData3 <= "0100100";
					SalidaData4 <= "0000010";
				when "0111111" => --63
					SalidaData3 <= "0110000";
					SalidaData4 <= "0000010";
				when "1000000" => --64
					SalidaData3 <= "0011001";
					SalidaData4 <= "0000010";
				when "1000001" => --65
					SalidaData3 <= "0010010";
					SalidaData4 <= "0000010";
				when "1000010" => --66
					SalidaData3 <= "0000010";
					SalidaData4 <= "0000010";
				when "1000011" => --67
					SalidaData3 <= "1111000";
					SalidaData4 <= "0000010";
				when "1000100" => --68
					SalidaData3 <= "0000000";
					SalidaData4 <= "0000010";
				when "1000101" => --69
					SalidaData3 <= "0010000";
					SalidaData4 <= "0000010";
				---- 70 al 79 ---------------
				when "1000110" => --70
					SalidaData3 <= "1000000";
					SalidaData4 <= "1111000";
				when "1000111" => --71
					SalidaData3 <= "1111001";
					SalidaData4 <= "1111000";
				when "1001000" => --72
					SalidaData3 <= "0100100";
					SalidaData4 <= "1111000";
				when "1001001" => --73
					SalidaData3 <= "0110000";
					SalidaData4 <= "1111000";
				when "1001010" => --74
					SalidaData3 <= "0011001";
					SalidaData4 <= "1111000";
				when "1001011" => --75
					SalidaData3 <= "0010010";
					SalidaData4 <= "1111000";
				when "1001100" => --76
					SalidaData3 <= "0000010";
					SalidaData4 <= "1111000";
				when "1001101" => --77
					SalidaData3 <= "1111000";
					SalidaData4 <= "1111000";
				when "1001110" => --78
					SalidaData3 <= "0000000";
					SalidaData4 <= "1111000";
				when "1001111" => --79
					SalidaData3 <= "0010000";
					SalidaData4 <= "1111000";
				---- 80 al 89 ---------------
				when "1010000" => --80
					SalidaData3 <= "1000000";
					SalidaData4 <= "0000000";
				when "1010001" => --81
					SalidaData3 <= "1111001";
					SalidaData4 <= "0000000";
				when "1010010" => --82
					SalidaData3 <= "0100100";
					SalidaData4 <= "0000000";
				when "1010011" => --83
					SalidaData3 <= "0110000";
					SalidaData4 <= "0000000";
				when "1010100" => --84
					SalidaData3 <= "0011001";
					SalidaData4 <= "0000000";
				when "1010101" => --85
					SalidaData3 <= "0010010";
					SalidaData4 <= "0000000";
				when "1010110" => --86
					SalidaData3 <= "0000010";
					SalidaData4 <= "0000000";
				when "1010111" => --87
					SalidaData3 <= "1111000";
					SalidaData4 <= "0000000";
				when "1011000" => --88
					SalidaData3 <= "0000000";
					SalidaData4 <= "0000000";
				when "1011001" => --89
					SalidaData3 <= "0010000";
					SalidaData4 <= "0000000";
				---- 80 al 89 ---------------
				when "1011010" => --90
					SalidaData3 <= "1000000";
					SalidaData4 <= "0010000";
				when "1011011" => --91
					SalidaData3 <= "1111001";
					SalidaData4 <= "0010000";
				when "1011100" => --92
					SalidaData3 <= "0100100";
					SalidaData4 <= "0010000";
				when "1011101" => --93
					SalidaData3 <= "0110000";
					SalidaData4 <= "0010000";
				when "1011110" => --94
					SalidaData3 <= "0011001";
					SalidaData4 <= "0010000";
				when "1011111" => --95
					SalidaData3 <= "0010010";
					SalidaData4 <= "0010000";
				when "1100000" => --96
					SalidaData3 <= "0000010";
					SalidaData4 <= "0010000";
				when "1100001" => --97
					SalidaData3 <= "1111000";
					SalidaData4 <= "0010000";
				when "1100010" => --98
					SalidaData3 <= "0000000";
					SalidaData4 <= "0010000";
				when "1100011" => --99
					SalidaData3 <= "0010000";
					SalidaData4 <= "0010000";
				when others =>
					SalidaData3 <= "1111111";
					SalidaData4 <= "1111111";
			end case;
		end process;
end architecture;