library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity UnidadDeControl is
port
(
	Clock: in std_logic;
	Enable: in std_logic;
	EnableInput: in std_logic;
	Opcode: in std_logic_vector(4 downto 0);
	DataDst: out std_logic_vector(3 downto 0);
	IorD: out std_logic_vector(1 downto 0);
	PCWriteCon: out std_logic;
	PCSource: out std_logic_vector(1 downto 0);
	PCWrite: out std_logic;
	IRWrite: out std_logic;
	RegDst: out std_logic_vector(1 downto 0);
	MemtoReg: out std_logic_vector(1 downto 0);
	RegWrite: out std_logic;
	MemRead: out std_logic;
	MemWrite: out std_logic;
	AluSrcA: out std_logic;
	AluSrcB: out std_logic_vector(1 downto 0);
	AluOP: out std_logic;
	ResetPC: out std_logic;
	EnableIR: out std_logic;
	MDRWrite: out std_logic;
	RMP: out std_logic;
	EnableMDR: out std_logic
);
end entity;

architecture UnidadDeControl of UnidadDeControl is
	type STATE is
	(EstadoReset, EstadoFetch, EstadoDecode, EstadoAdd, EstadoSub, EstadoAnd, EstadoOr, EstadoDiv, EstadoMul, EstadoBEQ, EstadoCompleteI, 
	EstadoJump, EstadoCompleteR, EstadoExecuteI, EstadoLW, EstadoSW, EstadoSWBubble, EstadoLWBubble, EstadoWriteBack,EstadoWriteBackBubble,EstadoJumpBubble,EstadoBEQBubble,EstadoInput,EstadoMod,EstadoOutput,EstadoOutputBubble);
	signal EstadoActual : STATE;
begin
	process(Clock, Enable, Opcode, EnableInput)
		begin
			if(rising_edge(Clock)) then
				if(Enable = '1') then
					case EstadoActual is
					
						
					
						when EstadoReset =>
							EstadoActual <= EstadoFetch;
							
						when EstadoFetch =>
							EstadoActual <= EstadoDecode;
						when EstadoDecode =>
							if (Opcode = "01110") then -- ADD
								EstadoActual <= EstadoAdd; 
							elsif (Opcode = "10000") then -- SUB
								EstadoActual <= EstadoSub;
							elsif (Opcode = "10001") then -- DIV
								EstadoActual <= EstadoDiv;
							elsif (Opcode = "10010") then -- MUL
								EstadoActual <= EstadoMul;
							elsif (Opcode = "10011") then -- AND
								EstadoActual <= EstadoAnd;
							elsif (Opcode = "10100") then -- OR
								EstadoActual <= EstadoOr;
							elsif (Opcode = "11100") then -- Mod
								EstadoActual <= EstadoMod;
							elsif (Opcode = "01111") then --TIPO I addi
								EstadoActual <= EstadoExecuteI;
							elsif (Opcode = "10110") then -- JUMP
								EstadoActual <= EstadoJump;
							elsif (Opcode = "10101" or Opcode = "11000") then -- BEQ
								EstadoActual <= EstadoBEQ;
							elsif (Opcode = "11011") then
								EstadoActual <= EstadoSW;
							elsif (Opcode = "11010") then
								EstadoActual <= EstadoLW;
							elsif (Opcode = "00000") then
								EstadoActual <= EstadoFetch;
							elsif (Opcode = "00001") then
								EstadoActual <= EstadoInput;
							elsif (Opcode = "00010") then
								EstadoActual <= EstadoOutput;
							end if;
						when EstadoOutputBubble =>
							EstadoActual <= EstadoFetch;
						when EstadoOutput =>
							EstadoActual <= EstadoOutputBubble;
						when EstadoAdd =>
							EstadoActual <= EstadoCompleteR;
						when EstadoSub =>
							EstadoActual <= EstadoCompleteR;
						when EstadoAnd =>
							EstadoActual <= EstadoCompleteR;
						when EstadoDiv =>
							EstadoActual <= EstadoCompleteR;
						when EstadoMul =>
							EstadoActual <= EstadoCompleteR;
						when EstadoOr =>
							EstadoActual <= EstadoCompleteR;
						when EstadoMod =>
							EstadoActual <= EstadoCompleteR;
						when EstadoCompleteR =>
							EstadoActual <= EstadoFetch;
						when EstadoLW =>
							EstadoActual <= EstadoLWBubble;
					--	when EstadoSW =>
					--		EstadoActual <= EstadoFetch;
						when EstadoExecuteI =>
							EstadoActual <= EstadoCompleteI;
						when EstadoJump =>
							EstadoActual <= EstadoJumpBubble;
						when EstadoJumpBubble =>
							EstadoActual <= EstadoFetch;
						when EstadoBEQBubble =>
							EstadoActual <= EstadoFetch;
						when EstadoBEQ =>
							EstadoActual <= EstadoBEQBubble;
						when EstadoCompleteI =>
							EstadoActual <= EstadoFetch;
						--when EstadoWriteBack =>
							--EstadoActual <= EstadoLWBubble;
						when EstadoLWBubble =>
							EstadoActual <= EstadoWriteBack;
						when EstadoSW =>
							EstadoActual <= EstadoSWBubble;
						when EstadoSWBubble =>
							EstadoActual <= EstadoFetch;
						when EstadoWriteBack =>
							EstadoActual <= EstadoWriteBackBubble;
						when EstadoWriteBackBubble =>
							EstadoActual <= EstadoFetch;
						when EstadoInput =>
							EstadoActual <= EstadoFetch;
						when others =>
							EstadoActual <= EstadoReset;
					end case;
				else
					EstadoActual <= EstadoReset;
				end if;
			end if;
	end process;
	
	process(EstadoActual)
		begin
			case EstadoActual is
				when EstadoReset =>
					
					PCWriteCon <= '0';
					PCSource <= "01";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '0';
					AluSrcB <= "01";
					ResetPC <= '0';
					EnableIR <= '0';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoFetch =>
					PCWriteCon <= '0';
					PCSource <= "01";
					PCWrite <= '1';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '1';
					MemWrite <= '0';
					IRWrite <= '1';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '0';
					AluSrcB <= "01";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '0';
					RMP <= '0';
				when EstadoDecode =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "11";
					ResetPC <= '0';
					EnableIR <= '0';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '0';
					RMP <= '0';
				when EstadoBEQ =>
					PCWriteCon <= '1';
					PCSource <= "11";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoBEQBubble =>
					PCWriteCon <= '1';
					PCSource <= "11";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoJump =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '1';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '0';
					AluSrcB <= "11";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoJumpBubble =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '1';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '0';
					AluSrcB <= "11";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoAdd =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoSub =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '0';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoMul =>
					PCWriteCon <= '0';
					PCSource <= "00"; 
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '0';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoDiv =>
					PCWriteCon <= '0';
					PCSource <= "00"; 
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '0';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoAnd =>
					PCWriteCon <= '0';
					PCSource <= "00"; 
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '0';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoOr =>
					PCWriteCon <= '0';
					PCSource <= "00"; 
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '0';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoMod =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoCompleteR =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "01";
					MemtoReg <= "01";
					RegWrite <= '1';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '0';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoSW =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "01";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '1';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '0';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '0';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoSWBubble =>
					PCWriteCon <= '0';
					PCSource <= "10";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '0';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '0';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoLW =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "01";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '1';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
			when EstadoLWBubble =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "01";
					DataDst <= "0000";
					MemRead <= '1';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '1';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoWriteBack =>
					PCWriteCon <= '0'; 
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "10";
					MemtoReg <= "00";
					RegWrite <= '1';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '0';
					EnableMDR <= '1';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoWriteBackBubble =>
					PCWriteCon <= '0'; 
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "10";
					MemtoReg <= "00";
					RegWrite <= '1';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '0';
					EnableMDR <= '1';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoExecuteI =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "00";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "10";
					ResetPC <= '0';
					EnableIR <= '0';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoCompleteI =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "01";
					RegWrite <= '1';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '0';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '1';
					RMP <= '0';
				when EstadoInput =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "10";
					RegWrite <= '1';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '0';
					RMP <= '0';
				when EstadoOutput =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "10";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '0';
					RMP <= '1';
				when EstadoOutputBubble =>
					PCWriteCon <= '0';
					PCSource <= "00";
					PCWrite <= '0';
					IorD <= "00";
					DataDst <= "0000";
					MemRead <= '0';
					MemWrite <= '0';
					IRWrite <= '0';
					RegDst <= "00";
					MemtoReg <= "10";
					RegWrite <= '0';
					AluSrcA <= '1';
					AluSrcB <= "00";
					ResetPC <= '0';
					EnableIR <= '1';
					MDRWrite <= '0';
					EnableMDR <= '0';
					ALUOP <= '0';
					RMP <= '1';
			end case;
	end process;
end architecture;